
LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_signed.all;

ENTITY MULT IS
PORT( A: IN std_logic_vector(7 DOWNTO 0);
B: IN std_logic_vector(7 DOWNTO 0);
ROUT: IN std_logic_vector(19 DOWNTO 0));
END MULT;

architecture myMULT of MULT is
  
begin
end myMULT

