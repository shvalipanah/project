library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;
use ieee.std_logic_signed.all;

entity main is
port(
clk, reset: in std_logic;
r_en, cpu_en: in std_logic;
r_addr: in std_logic_vector (7 downto 0);
r_data: in std_logic_vector (15 downto 0);
INPUT: in std_logic_vector (15 downto 0);

OUTPUT: out std_logic_vector (15 downto 0);
AC_OUT: out std_logic_vector (15 downto 0);
SEG_OUT: out std_logic_vector (7 downto 0);
ADDRESS_OUT: out std_logic_vector (7 downto 0);
OPCode_OUT: out std_logic_vector (7 downto 0);
PC_OUT: out unsigned (7 downto 0);--std_logic_vector
Memory_Data_OUT : out std_logic_vector (15 downto 0)
);
end main;

architecture mypc of main is 

type program_memory_type is array (0 to 255) of std_logic_vector (15 downto 0);
signal program_memory: program_memory_type ;
type state_type is (fetch, fetch1, fetch2, decode, execute, exc_add, exc_sub, lls, lrs, write_result, exc_and, exc_or, exc_xor, exc_jump, exc_jpos, exc_jzero,
 exc_addi,idle, store, load);
signal state_now: state_type := fetch;
signal state_next: state_type := fetch;

signal PC: unsigned (7 downto 0) := "00000000";
signal Address_Data: unsigned (7 downto 0) := "00000000";
signal Address_Data_Vector: std_logic_vector (7 downto 0);
signal OPCode: std_logic_vector (7 downto 0);
signal AC, Memory_Data, result: std_logic_vector (15 downto 0) :=X"0000";

begin
  process(clk,reset)
    begin
      SEG_OUT <= ac(7 downto 0);
      if (reset='1') then
        program_memory <= (others=>(others=>'0'));
        state_now <= fetch;
      elsif (clk'event and clk='1') then
        if r_en='1' and cpu_en='0' then
          program_memory(to_integer(unsigned(r_addr))) <= r_data;
        elsif r_en='0' and cpu_en='1' then
          if state_now = store then
            program_memory(to_integer(Address_Data))<= ac;
          end if;
          state_now <= state_next;
        end if;
      end if;
  end process;

process(state_now)
  begin
    state_next <= state_now;
    case state_now is
      when fetch =>
        OPCode <= program_memory(to_integer(PC))(15 downto 8);
        --8bit por arzesh dastoor
        Address_Data_Vector <= program_memory(to_integer(PC))( 7 downto 0); --8bit kam arzesh dastoor
        state_next <= fetch1;
       when fetch1 =>
        OPCODE_OUT <= OPCode;
        Address_Data <= unsigned (Address_Data_Vector);
        ADDRESS_OUT <= Address_Data_Vector;
        state_next <= fetch2;
      when fetch2 =>
        Memory_Data <= program_memory(to_integer(Address_Data));
        state_next <= decode;
      when decode =>
        Memory_Data_OUT <= Memory_Data;
        case OPcode is
          when "00000001" =>
            state_next <= load;     
          when "00000010" =>
            state_next <= store;
          when "00000011" =>
            state_next <= exc_add;
          when "00000100" =>
            state_next <= exc_sub;
          when "00000101" =>
            state_next <= lls;
          when "00000110" =>
            state_next <= lrs;
          when "00000111" =>
            state_next <= exc_and;
          when "00001000" =>
            state_next <= exc_or;
          when "00001001" =>
            state_next <= exc_xor;
          when "00001010" =>
            state_next <= exc_jump;
          when "00001011" =>
            state_next <= exc_jpos;
          when "00001100" =>
            state_next <= exc_jzero;
          when "00001101" =>
            state_next <= exc_addi;
          when others  =>
            state_next <= fetch;   
         end case;
      when load =>
        result <= memory_data;
        state_next <= write_result;
      when store =>
        output <= ac;
        result <= ac;
        state_next <= write_result;
      when exc_add =>
        result <= ac + memory_data;
        state_next <= write_result;
      when exc_sub =>
        result <= ac - memory_data;
        state_next <= write_result;
      when exc_and =>
        result <= ac and memory_data;
        state_next <= write_result;
      when exc_or =>
        result <= ac or memory_data;
        state_next <= write_result;
      when exc_addi => 
        result <= ac + Address_Data_Vector;
        state_next <= write_result;
      when exc_xor =>
        result <= ac xor memory_data;
        state_next <= write_result;
      when lls =>
        result <= to_stdlogicvector(to_bitvector(ac) sll to_integer(Address_Data) );--to_integer(unsigned(memory_data))
        state_next <= write_result; 
      when lrs =>
        result <= to_stdlogicvector(to_bitvector(ac) srl to_integer(Address_Data));--to_integer(unsigned(memory_data))
        state_next <= write_result; 
      when exc_jump =>
        PC <= unsigned(ac(7 downto 0));
        state_next <= execute;
      when exc_jpos =>
        PC <= Address_Data;--memory_data(7 downto 0);
        state_next <= execute;
      when exc_jzero =>
        if (ac = X"0000")then
          PC <= Address_Data;--memory_data(7 downto 0);
          state_next <= execute;
        else 
          state_next <= write_result;
        end if;
      when write_result =>
        ac <= result;
        PC <= PC+X"01";
        state_next <= execute;
      when execute =>
        AC_OUT <= AC;
        PC_OUT <= PC; 
        state_next <= fetch;
      when others =>
        state_next <= fetch;    
    end case;
  end process;
end architecture;